LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY Regn IS
PORT (
	RST, CLK : IN STD_LOGIC;
	En : IN STD_LOGIC;
	D : IN INTEGER;
	Q : OUT INTEGER
);
END Regn;

ARCHITECTURE RTL OF Regn IS
BEGIN
PROCESS (RST, CLK)
BEGIN
IF (RST = '1') THEN
	Q <= 0;
ELSIF (CLK'EVENT and CLK = '1') THEN 
	IF (EN = '1') THEN
		Q <= D;
	END IF;
END IF;
END PROCESS;

END RTL; 